`timescale 1ns/1ps

// latency = 4

// Fully pipeline PINI circuit in 4 clock cycles.
// This file has been automatically generated.
`ifdef FULLVERIF
(* fv_prop = "PINI", fv_strat = "composite", fv_order=d *)
`endif
module bp_c_common # ( parameter d=2 ) (
    clk,
    t1,
    t2,
    t3,
    t4,
    t5,
    t6,
    t7,
    t8,
    t9,
    t10,
    t11,
    t12,
    t13,
    t14,
    t15,
    t16,
    t17,
    t18,
    t19,
    t20,
    t21,
    t22,
    t23,
    t24,
    t25,
    t26,
    t27,
    ds,
    m1,
    m2,
    m3,
    m4,
    m5,
    m6,
    m7,
    m8,
    m9,
    m10,
    m11,
    m12,
    m13,
    m14,
    m15,
    m16,
    m17,
    m18,
    m19,
    m20,
    m21,
    m22,
    m23,
    m24,
    m25,
    m26,
    m27,
    m28,
    m29,
    m30,
    m31,
    m32,
    m33,
    m34,
    m35,
    m36,
    m37,
    m38,
    m39,
    m40,
    m41,
    m42,
    m43,
    m44,
    m45,
    m46,
    m47,
    m48,
    m49,
    m50,
    m51,
    m52,
    m53,
    m54,
    m55,
    m56,
    m57,
    m58,
    m59,
    m60,
    m61,
    m62,
    m63,
    rnd_0,
    rnd_1,
    rnd_2,
);
`include "MSKand_hpc1.vh"
`include "MSKand_hpc2.vh"
`include "MSKand_hpc3.vh"
(* fv_type="clock" *)
input clk;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t1;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t2;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t3;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t4;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t5;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t6;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t7;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t8;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t9;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t10;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t11;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t12;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t13;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t14;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t15;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t16;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t17;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t18;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t19;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t20;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t21;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t22;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t23;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t24;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t25;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t26;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] t27;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] ds;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m1;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m2;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m3;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m4;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m5;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m6;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m7;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m8;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m9;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m10;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m11;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m12;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m13;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m14;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m15;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m16;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m17;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m18;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m19;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m20;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m21;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m22;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m23;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m24;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m25;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m26;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m27;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m28;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m29;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m30;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m31;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m32;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m33;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m34;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m35;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m36;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m37;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m38;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m39;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m40;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m41;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m42;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m43;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m44;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m45;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m46;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m47;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m48;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m49;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m50;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m51;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m52;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m53;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m54;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m55;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m56;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m57;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m58;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m59;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m60;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m61;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m62;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] m63;
(* fv_type="random", fv_count=1, fv_rnd_count_0=9*(1*d*(d-1)), fv_rnd_lat_0=0  *)
input [9*(1*d*(d-1))-1:0] rnd_0;
(* fv_type="random", fv_count=1, fv_rnd_count_0=3*(1*d*(d-1))+4*(1*d*(d-1)/2), fv_rnd_lat_0=1  *)
input [3*(1*d*(d-1))+4*(1*d*(d-1)/2)-1:0] rnd_1;
(* fv_type="random", fv_count=1, fv_rnd_count_0=18*(1*d*(d-1)/2), fv_rnd_lat_0=2  *)
input [18*(1*d*(d-1)/2)-1:0] rnd_2;
wire [d-1:0] ds_0;
wire [d-1:0] ds_1;
wire [d-1:0] ds_2;
wire [d-1:0] ds_3;
wire [d-1:0] m1_1;
wire [d-1:0] m1_2;
wire [d-1:0] m1_3;
wire [d-1:0] m1_4;
wire [d-1:0] m10_1;
wire [d-1:0] m10_2;
wire [d-1:0] m10_3;
wire [d-1:0] m10_4;
wire [d-1:0] m11_1;
wire [d-1:0] m11_2;
wire [d-1:0] m11_3;
wire [d-1:0] m11_4;
wire [d-1:0] m12_1;
wire [d-1:0] m12_2;
wire [d-1:0] m12_3;
wire [d-1:0] m12_4;
wire [d-1:0] m13_1;
wire [d-1:0] m13_2;
wire [d-1:0] m13_3;
wire [d-1:0] m13_4;
wire [d-1:0] m14_1;
wire [d-1:0] m14_2;
wire [d-1:0] m14_3;
wire [d-1:0] m14_4;
wire [d-1:0] m15_1;
wire [d-1:0] m15_2;
wire [d-1:0] m15_3;
wire [d-1:0] m15_4;
wire [d-1:0] m16_1;
wire [d-1:0] m16_2;
wire [d-1:0] m16_3;
wire [d-1:0] m16_4;
wire [d-1:0] m17_1;
wire [d-1:0] m17_2;
wire [d-1:0] m17_3;
wire [d-1:0] m17_4;
wire [d-1:0] m18_1;
wire [d-1:0] m18_2;
wire [d-1:0] m18_3;
wire [d-1:0] m18_4;
wire [d-1:0] m19_1;
wire [d-1:0] m19_2;
wire [d-1:0] m19_3;
wire [d-1:0] m19_4;
wire [d-1:0] m2_1;
wire [d-1:0] m2_2;
wire [d-1:0] m2_3;
wire [d-1:0] m2_4;
wire [d-1:0] m20_1;
wire [d-1:0] m20_2;
wire [d-1:0] m20_3;
wire [d-1:0] m20_4;
wire [d-1:0] m21_1;
wire [d-1:0] m21_2;
wire [d-1:0] m21_3;
wire [d-1:0] m21_4;
wire [d-1:0] m22_1;
wire [d-1:0] m22_2;
wire [d-1:0] m22_3;
wire [d-1:0] m22_4;
wire [d-1:0] m23_1;
wire [d-1:0] m23_2;
wire [d-1:0] m23_3;
wire [d-1:0] m23_4;
wire [d-1:0] m24_1;
wire [d-1:0] m24_2;
wire [d-1:0] m24_3;
wire [d-1:0] m24_4;
wire [d-1:0] m25_2;
wire [d-1:0] m25_3;
wire [d-1:0] m25_4;
wire [d-1:0] m26_2;
wire [d-1:0] m26_3;
wire [d-1:0] m26_4;
wire [d-1:0] m27_1;
wire [d-1:0] m27_2;
wire [d-1:0] m27_3;
wire [d-1:0] m27_4;
wire [d-1:0] m28_2;
wire [d-1:0] m28_3;
wire [d-1:0] m28_4;
wire [d-1:0] m29_3;
wire [d-1:0] m29_4;
wire [d-1:0] m3_1;
wire [d-1:0] m3_2;
wire [d-1:0] m3_3;
wire [d-1:0] m3_4;
wire [d-1:0] m30_3;
wire [d-1:0] m30_4;
wire [d-1:0] m31_2;
wire [d-1:0] m31_3;
wire [d-1:0] m31_4;
wire [d-1:0] m32_3;
wire [d-1:0] m32_4;
wire [d-1:0] m33_3;
wire [d-1:0] m33_4;
wire [d-1:0] m34_2;
wire [d-1:0] m34_3;
wire [d-1:0] m34_4;
wire [d-1:0] m35_3;
wire [d-1:0] m35_4;
wire [d-1:0] m36_3;
wire [d-1:0] m36_4;
wire [d-1:0] m37_3;
wire [d-1:0] m37_4;
wire [d-1:0] m38_3;
wire [d-1:0] m38_4;
wire [d-1:0] m39_3;
wire [d-1:0] m39_4;
wire [d-1:0] m4_1;
wire [d-1:0] m4_2;
wire [d-1:0] m4_3;
wire [d-1:0] m4_4;
wire [d-1:0] m40_3;
wire [d-1:0] m40_4;
wire [d-1:0] m41_3;
wire [d-1:0] m41_4;
wire [d-1:0] m42_3;
wire [d-1:0] m42_4;
wire [d-1:0] m43_3;
wire [d-1:0] m43_4;
wire [d-1:0] m44_3;
wire [d-1:0] m44_4;
wire [d-1:0] m45_3;
wire [d-1:0] m45_4;
wire [d-1:0] m46_4;
wire [d-1:0] m47_4;
wire [d-1:0] m48_4;
wire [d-1:0] m49_4;
wire [d-1:0] m5_1;
wire [d-1:0] m5_2;
wire [d-1:0] m5_3;
wire [d-1:0] m5_4;
wire [d-1:0] m50_4;
wire [d-1:0] m51_4;
wire [d-1:0] m52_4;
wire [d-1:0] m53_4;
wire [d-1:0] m54_4;
wire [d-1:0] m55_4;
wire [d-1:0] m56_4;
wire [d-1:0] m57_4;
wire [d-1:0] m58_4;
wire [d-1:0] m59_4;
wire [d-1:0] m6_1;
wire [d-1:0] m6_2;
wire [d-1:0] m6_3;
wire [d-1:0] m6_4;
wire [d-1:0] m60_4;
wire [d-1:0] m61_4;
wire [d-1:0] m62_4;
wire [d-1:0] m63_4;
wire [d-1:0] m7_1;
wire [d-1:0] m7_2;
wire [d-1:0] m7_3;
wire [d-1:0] m7_4;
wire [d-1:0] m8_1;
wire [d-1:0] m8_2;
wire [d-1:0] m8_3;
wire [d-1:0] m8_4;
wire [d-1:0] m9_1;
wire [d-1:0] m9_2;
wire [d-1:0] m9_3;
wire [d-1:0] m9_4;
wire [d-1:0] t1_0;
wire [d-1:0] t1_1;
wire [d-1:0] t1_2;
wire [d-1:0] t1_3;
wire [d-1:0] t10_0;
wire [d-1:0] t10_1;
wire [d-1:0] t10_2;
wire [d-1:0] t10_3;
wire [d-1:0] t11_0;
wire [d-1:0] t12_0;
wire [d-1:0] t13_0;
wire [d-1:0] t13_1;
wire [d-1:0] t13_2;
wire [d-1:0] t13_3;
wire [d-1:0] t14_0;
wire [d-1:0] t14_1;
wire [d-1:0] t15_0;
wire [d-1:0] t15_1;
wire [d-1:0] t15_2;
wire [d-1:0] t15_3;
wire [d-1:0] t16_0;
wire [d-1:0] t16_1;
wire [d-1:0] t16_2;
wire [d-1:0] t16_3;
wire [d-1:0] t17_0;
wire [d-1:0] t17_1;
wire [d-1:0] t17_2;
wire [d-1:0] t17_3;
wire [d-1:0] t18_0;
wire [d-1:0] t19_0;
wire [d-1:0] t19_1;
wire [d-1:0] t19_2;
wire [d-1:0] t19_3;
wire [d-1:0] t2_0;
wire [d-1:0] t2_1;
wire [d-1:0] t2_2;
wire [d-1:0] t2_3;
wire [d-1:0] t20_0;
wire [d-1:0] t20_1;
wire [d-1:0] t20_2;
wire [d-1:0] t20_3;
wire [d-1:0] t21_0;
wire [d-1:0] t22_0;
wire [d-1:0] t22_1;
wire [d-1:0] t22_2;
wire [d-1:0] t22_3;
wire [d-1:0] t23_0;
wire [d-1:0] t23_1;
wire [d-1:0] t23_2;
wire [d-1:0] t23_3;
wire [d-1:0] t24_0;
wire [d-1:0] t24_1;
wire [d-1:0] t25_0;
wire [d-1:0] t25_1;
wire [d-1:0] t26_0;
wire [d-1:0] t26_1;
wire [d-1:0] t27_0;
wire [d-1:0] t27_1;
wire [d-1:0] t27_2;
wire [d-1:0] t27_3;
wire [d-1:0] t3_0;
wire [d-1:0] t3_1;
wire [d-1:0] t3_2;
wire [d-1:0] t3_3;
wire [d-1:0] t4_0;
wire [d-1:0] t4_1;
wire [d-1:0] t4_2;
wire [d-1:0] t4_3;
wire [d-1:0] t5_0;
wire [d-1:0] t6_0;
wire [d-1:0] t6_1;
wire [d-1:0] t6_2;
wire [d-1:0] t6_3;
wire [d-1:0] t7_0;
wire [d-1:0] t8_0;
wire [d-1:0] t8_1;
wire [d-1:0] t8_2;
wire [d-1:0] t8_3;
wire [d-1:0] t9_0;
wire [d-1:0] t9_1;
wire [d-1:0] t9_2;
wire [d-1:0] t9_3;
assign t1_0 = t1;
assign t2_0 = t2;
assign t3_0 = t3;
assign t4_0 = t4;
assign t5_0 = t5;
assign t6_0 = t6;
assign t7_0 = t7;
assign t8_0 = t8;
assign t9_0 = t9;
assign t10_0 = t10;
assign t11_0 = t11;
assign t12_0 = t12;
assign t13_0 = t13;
assign t14_0 = t14;
assign t15_0 = t15;
assign t16_0 = t16;
assign t17_0 = t17;
assign t18_0 = t18;
assign t19_0 = t19;
assign t20_0 = t20;
assign t21_0 = t21;
assign t22_0 = t22;
assign t23_0 = t23;
assign t24_0 = t24;
assign t25_0 = t25;
assign t26_0 = t26;
assign t27_0 = t27;
assign ds_0 = ds;
assign m1 = m1_4;
assign m2 = m2_4;
assign m3 = m3_4;
assign m4 = m4_4;
assign m5 = m5_4;
assign m6 = m6_4;
assign m7 = m7_4;
assign m8 = m8_4;
assign m9 = m9_4;
assign m10 = m10_4;
assign m11 = m11_4;
assign m12 = m12_4;
assign m13 = m13_4;
assign m14 = m14_4;
assign m15 = m15_4;
assign m16 = m16_4;
assign m17 = m17_4;
assign m18 = m18_4;
assign m19 = m19_4;
assign m20 = m20_4;
assign m21 = m21_4;
assign m22 = m22_4;
assign m23 = m23_4;
assign m24 = m24_4;
assign m25 = m25_4;
assign m26 = m26_4;
assign m27 = m27_4;
assign m28 = m28_4;
assign m29 = m29_4;
assign m30 = m30_4;
assign m31 = m31_4;
assign m32 = m32_4;
assign m33 = m33_4;
assign m34 = m34_4;
assign m35 = m35_4;
assign m36 = m36_4;
assign m37 = m37_4;
assign m38 = m38_4;
assign m39 = m39_4;
assign m40 = m40_4;
assign m41 = m41_4;
assign m42 = m42_4;
assign m43 = m43_4;
assign m44 = m44_4;
assign m45 = m45_4;
assign m46 = m46_4;
assign m47 = m47_4;
assign m48 = m48_4;
assign m49 = m49_4;
assign m50 = m50_4;
assign m51 = m51_4;
assign m52 = m52_4;
assign m53 = m53_4;
assign m54 = m54_4;
assign m55 = m55_4;
assign m56 = m56_4;
assign m57 = m57_4;
assign m58 = m58_4;
assign m59 = m59_4;
assign m60 = m60_4;
assign m61 = m61_4;
assign m62 = m62_4;
assign m63 = m63_4;




MSKand_hpc3o #(.d(d)) comp_m1_1 (
    .out(m1_1),
    .rnd(rnd_0[0 +: 1*d*(d-1)]),
    .ina(t13_0),
    .ina_prev(t13_1),
    .inb(t6_0),
    .clk(clk)
);
MSKand_hpc3o_swapped #(.d(d)) comp_m2_1 (
    .out(m2_1),
    .rnd(rnd_0[1*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t23_0),
    .inb(t8_0),
    .inb_prev(t8_1),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m3_1 (
    .out(m3_1),
    .ina(t14_1),
    .inb(m1_1)
);
MSKand_hpc3o_swapped #(.d(d)) comp_m4_1 (
    .out(m4_1),
    .rnd(rnd_0[2*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t19_0),
    .inb(ds_0),
    .inb_prev(ds_1),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m5_1 (
    .out(m5_1),
    .ina(m4_1),
    .inb(m1_1)
);
MSKand_hpc3o #(.d(d)) comp_m6_1 (
    .out(m6_1),
    .rnd(rnd_0[3*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t3_0),
    .ina_prev(t3_1),
    .inb(t16_0),
    .clk(clk)
);
MSKand_hpc3o #(.d(d)) comp_m7_1 (
    .out(m7_1),
    .rnd(rnd_0[4*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t22_0),
    .ina_prev(t22_1),
    .inb(t9_0),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m8_1 (
    .out(m8_1),
    .ina(t26_1),
    .inb(m6_1)
);
MSKand_hpc3o #(.d(d)) comp_m9_1 (
    .out(m9_1),
    .rnd(rnd_0[5*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t20_0),
    .ina_prev(t20_1),
    .inb(t17_0),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m10_1 (
    .out(m10_1),
    .ina(m9_1),
    .inb(m6_1)
);
MSKand_hpc3o #(.d(d)) comp_m11_1 (
    .out(m11_1),
    .rnd(rnd_0[6*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t1_0),
    .ina_prev(t1_1),
    .inb(t15_0),
    .clk(clk)
);
MSKand_hpc3o_swapped #(.d(d)) comp_m12_1 (
    .out(m12_1),
    .rnd(rnd_0[7*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t4_0),
    .inb(t27_0),
    .inb_prev(t27_1),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m13_1 (
    .out(m13_1),
    .ina(m12_1),
    .inb(m11_1)
);
MSKand_hpc3o #(.d(d)) comp_m14_1 (
    .out(m14_1),
    .rnd(rnd_0[8*(1*d*(d-1)) +: 1*d*(d-1)]),
    .ina(t2_0),
    .ina_prev(t2_1),
    .inb(t10_0),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m15_1 (
    .out(m15_1),
    .ina(m14_1),
    .inb(m11_1)
);
MSKxor #(.d(d)) comp_m16_1 (
    .out(m16_1),
    .ina(m3_1),
    .inb(m2_1)
);
MSKxor #(.d(d)) comp_m17_1 (
    .out(m17_1),
    .ina(m5_1),
    .inb(t24_1)
);
MSKxor #(.d(d)) comp_m18_1 (
    .out(m18_1),
    .ina(m8_1),
    .inb(m7_1)
);
MSKxor #(.d(d)) comp_m19_1 (
    .out(m19_1),
    .ina(m10_1),
    .inb(m15_1)
);
MSKxor #(.d(d)) comp_m20_1 (
    .out(m20_1),
    .ina(m16_1),
    .inb(m13_1)
);
MSKxor #(.d(d)) comp_m21_1 (
    .out(m21_1),
    .ina(m17_1),
    .inb(m15_1)
);
MSKxor #(.d(d)) comp_m22_1 (
    .out(m22_1),
    .ina(m18_1),
    .inb(m13_1)
);
MSKxor #(.d(d)) comp_m23_1 (
    .out(m23_1),
    .ina(m19_1),
    .inb(t25_1)
);
MSKxor #(.d(d)) comp_m24_1 (
    .out(m24_1),
    .ina(m22_1),
    .inb(m23_1)
);
MSKand_hpc3o #(.d(d)) comp_m25_2 (
    .out(m25_2),
    .rnd(rnd_1[0 +: 1*d*(d-1)]),
    .ina(m22_1),
    .ina_prev(m22_2),
    .inb(m20_1),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m26_2 (
    .out(m26_2),
    .ina(m21_2),
    .inb(m25_2)
);
MSKxor #(.d(d)) comp_m27_1 (
    .out(m27_1),
    .ina(m20_1),
    .inb(m21_1)
);
MSKxor #(.d(d)) comp_m28_2 (
    .out(m28_2),
    .ina(m23_2),
    .inb(m25_2)
);
MSKand_hpc2o #(.d(d)) comp_m29_3 (
    .out(m29_3),
    .rnd(rnd_1[1*(1*d*(d-1)) +: 1*d*(d-1)/2]),
    .ina(m28_2),
    .inb(m27_1),
    .inb_prev(m27_2),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m30_3 (
    .out(m30_3),
    .rnd(rnd_1[1*(1*d*(d-1))+1*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m26_2),
    .inb(m24_1),
    .inb_prev(m24_2),
    .clk(clk)
);
MSKand_hpc3o_swapped #(.d(d)) comp_m31_2 (
    .out(m31_2),
    .rnd(rnd_1[1*(1*d*(d-1))+2*(1*d*(d-1)/2) +: 1*d*(d-1)]),
    .ina(m20_1),
    .inb(m23_1),
    .inb_prev(m23_2),
    .clk(clk)
);
MSKand_hpc2o_swapped #(.d(d)) comp_m32_3 (
    .out(m32_3),
    .rnd(rnd_1[2*(1*d*(d-1))+2*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m27_1),
    .ina_prev(m27_2),
    .inb(m31_2),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m33_3 (
    .out(m33_3),
    .ina(m27_3),
    .inb(m25_3)
);
MSKand_hpc3o #(.d(d)) comp_m34_2 (
    .out(m34_2),
    .rnd(rnd_1[2*(1*d*(d-1))+3*(1*d*(d-1)/2) +: 1*d*(d-1)]),
    .ina(m21_1),
    .ina_prev(m21_2),
    .inb(m22_1),
    .clk(clk)
);
MSKand_hpc2o_swapped #(.d(d)) comp_m35_3 (
    .out(m35_3),
    .rnd(rnd_1[3*(1*d*(d-1))+3*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m24_1),
    .ina_prev(m24_2),
    .inb(m34_2),
    .clk(clk)
);
MSKxor #(.d(d)) comp_m36_3 (
    .out(m36_3),
    .ina(m24_3),
    .inb(m25_3)
);
MSKxor #(.d(d)) comp_m37_3 (
    .out(m37_3),
    .ina(m21_3),
    .inb(m29_3)
);
MSKxor #(.d(d)) comp_m38_3 (
    .out(m38_3),
    .ina(m32_3),
    .inb(m33_3)
);
MSKxor #(.d(d)) comp_m39_3 (
    .out(m39_3),
    .ina(m23_3),
    .inb(m30_3)
);
MSKxor #(.d(d)) comp_m40_3 (
    .out(m40_3),
    .ina(m35_3),
    .inb(m36_3)
);
MSKxor #(.d(d)) comp_m41_3 (
    .out(m41_3),
    .ina(m38_3),
    .inb(m40_3)
);
MSKxor #(.d(d)) comp_m42_3 (
    .out(m42_3),
    .ina(m37_3),
    .inb(m39_3)
);
MSKxor #(.d(d)) comp_m43_3 (
    .out(m43_3),
    .ina(m37_3),
    .inb(m38_3)
);
MSKxor #(.d(d)) comp_m44_3 (
    .out(m44_3),
    .ina(m39_3),
    .inb(m40_3)
);
MSKxor #(.d(d)) comp_m45_3 (
    .out(m45_3),
    .ina(m42_3),
    .inb(m41_3)
);
MSKand_hpc2o #(.d(d)) comp_m46_4 (
    .out(m46_4),
    .rnd(rnd_2[0 +: 1*d*(d-1)/2]),
    .ina(m44_3),
    .inb(t6_2),
    .inb_prev(t6_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m47_4 (
    .out(m47_4),
    .rnd(rnd_2[1*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m40_3),
    .inb(t8_2),
    .inb_prev(t8_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m48_4 (
    .out(m48_4),
    .rnd(rnd_2[2*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m39_3),
    .inb(ds_2),
    .inb_prev(ds_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m49_4 (
    .out(m49_4),
    .rnd(rnd_2[3*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m43_3),
    .inb(t16_2),
    .inb_prev(t16_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m50_4 (
    .out(m50_4),
    .rnd(rnd_2[4*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m38_3),
    .inb(t9_2),
    .inb_prev(t9_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m51_4 (
    .out(m51_4),
    .rnd(rnd_2[5*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m37_3),
    .inb(t17_2),
    .inb_prev(t17_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m52_4 (
    .out(m52_4),
    .rnd(rnd_2[6*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m42_3),
    .inb(t15_2),
    .inb_prev(t15_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m53_4 (
    .out(m53_4),
    .rnd(rnd_2[7*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m45_3),
    .inb(t27_2),
    .inb_prev(t27_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m54_4 (
    .out(m54_4),
    .rnd(rnd_2[8*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m41_3),
    .inb(t10_2),
    .inb_prev(t10_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m55_4 (
    .out(m55_4),
    .rnd(rnd_2[9*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m44_3),
    .inb(t13_2),
    .inb_prev(t13_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m56_4 (
    .out(m56_4),
    .rnd(rnd_2[10*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m40_3),
    .inb(t23_2),
    .inb_prev(t23_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m57_4 (
    .out(m57_4),
    .rnd(rnd_2[11*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m39_3),
    .inb(t19_2),
    .inb_prev(t19_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m58_4 (
    .out(m58_4),
    .rnd(rnd_2[12*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m43_3),
    .inb(t3_2),
    .inb_prev(t3_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m59_4 (
    .out(m59_4),
    .rnd(rnd_2[13*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m38_3),
    .inb(t22_2),
    .inb_prev(t22_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m60_4 (
    .out(m60_4),
    .rnd(rnd_2[14*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m37_3),
    .inb(t20_2),
    .inb_prev(t20_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m61_4 (
    .out(m61_4),
    .rnd(rnd_2[15*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m42_3),
    .inb(t1_2),
    .inb_prev(t1_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m62_4 (
    .out(m62_4),
    .rnd(rnd_2[16*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m45_3),
    .inb(t4_2),
    .inb_prev(t4_3),
    .clk(clk)
);
MSKand_hpc2o #(.d(d)) comp_m63_4 (
    .out(m63_4),
    .rnd(rnd_2[17*(1*d*(d-1)/2) +: 1*d*(d-1)/2]),
    .ina(m41_3),
    .inb(t2_2),
    .inb_prev(t2_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m4_1 (
    .in(m4_1),
    .out(m4_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m4_2 (
    .in(m4_2),
    .out(m4_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m4_3 (
    .in(m4_3),
    .out(m4_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m30_3 (
    .in(m30_3),
    .out(m30_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m18_1 (
    .in(m18_1),
    .out(m18_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m18_2 (
    .in(m18_2),
    .out(m18_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m18_3 (
    .in(m18_3),
    .out(m18_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t9_0 (
    .in(t9_0),
    .out(t9_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t9_1 (
    .in(t9_1),
    .out(t9_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t9_2 (
    .in(t9_2),
    .out(t9_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t3_0 (
    .in(t3_0),
    .out(t3_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t3_1 (
    .in(t3_1),
    .out(t3_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t3_2 (
    .in(t3_2),
    .out(t3_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t6_0 (
    .in(t6_0),
    .out(t6_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t6_1 (
    .in(t6_1),
    .out(t6_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t6_2 (
    .in(t6_2),
    .out(t6_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m40_3 (
    .in(m40_3),
    .out(m40_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t19_0 (
    .in(t19_0),
    .out(t19_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t19_1 (
    .in(t19_1),
    .out(t19_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t19_2 (
    .in(t19_2),
    .out(t19_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t14_0 (
    .in(t14_0),
    .out(t14_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m13_1 (
    .in(m13_1),
    .out(m13_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m13_2 (
    .in(m13_2),
    .out(m13_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m13_3 (
    .in(m13_3),
    .out(m13_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m7_1 (
    .in(m7_1),
    .out(m7_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m7_2 (
    .in(m7_2),
    .out(m7_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m7_3 (
    .in(m7_3),
    .out(m7_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m32_3 (
    .in(m32_3),
    .out(m32_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m10_1 (
    .in(m10_1),
    .out(m10_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m10_2 (
    .in(m10_2),
    .out(m10_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m10_3 (
    .in(m10_3),
    .out(m10_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m12_1 (
    .in(m12_1),
    .out(m12_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m12_2 (
    .in(m12_2),
    .out(m12_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m12_3 (
    .in(m12_3),
    .out(m12_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m23_1 (
    .in(m23_1),
    .out(m23_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m23_2 (
    .in(m23_2),
    .out(m23_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m23_3 (
    .in(m23_3),
    .out(m23_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m31_2 (
    .in(m31_2),
    .out(m31_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m31_3 (
    .in(m31_3),
    .out(m31_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_ds_0 (
    .in(ds_0),
    .out(ds_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_ds_1 (
    .in(ds_1),
    .out(ds_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_ds_2 (
    .in(ds_2),
    .out(ds_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m34_2 (
    .in(m34_2),
    .out(m34_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m34_3 (
    .in(m34_3),
    .out(m34_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t8_0 (
    .in(t8_0),
    .out(t8_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t8_1 (
    .in(t8_1),
    .out(t8_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t8_2 (
    .in(t8_2),
    .out(t8_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m26_2 (
    .in(m26_2),
    .out(m26_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m26_3 (
    .in(m26_3),
    .out(m26_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t20_0 (
    .in(t20_0),
    .out(t20_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t20_1 (
    .in(t20_1),
    .out(t20_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t20_2 (
    .in(t20_2),
    .out(t20_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m20_1 (
    .in(m20_1),
    .out(m20_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m20_2 (
    .in(m20_2),
    .out(m20_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m20_3 (
    .in(m20_3),
    .out(m20_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m36_3 (
    .in(m36_3),
    .out(m36_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m29_3 (
    .in(m29_3),
    .out(m29_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t27_0 (
    .in(t27_0),
    .out(t27_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t27_1 (
    .in(t27_1),
    .out(t27_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t27_2 (
    .in(t27_2),
    .out(t27_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t23_0 (
    .in(t23_0),
    .out(t23_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t23_1 (
    .in(t23_1),
    .out(t23_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t23_2 (
    .in(t23_2),
    .out(t23_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m16_1 (
    .in(m16_1),
    .out(m16_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m16_2 (
    .in(m16_2),
    .out(m16_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m16_3 (
    .in(m16_3),
    .out(m16_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t13_0 (
    .in(t13_0),
    .out(t13_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t13_1 (
    .in(t13_1),
    .out(t13_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t13_2 (
    .in(t13_2),
    .out(t13_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t26_0 (
    .in(t26_0),
    .out(t26_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m37_3 (
    .in(m37_3),
    .out(m37_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m3_1 (
    .in(m3_1),
    .out(m3_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m3_2 (
    .in(m3_2),
    .out(m3_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m3_3 (
    .in(m3_3),
    .out(m3_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m17_1 (
    .in(m17_1),
    .out(m17_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m17_2 (
    .in(m17_2),
    .out(m17_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m17_3 (
    .in(m17_3),
    .out(m17_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m39_3 (
    .in(m39_3),
    .out(m39_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m22_1 (
    .in(m22_1),
    .out(m22_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m22_2 (
    .in(m22_2),
    .out(m22_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m22_3 (
    .in(m22_3),
    .out(m22_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m2_1 (
    .in(m2_1),
    .out(m2_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m2_2 (
    .in(m2_2),
    .out(m2_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m2_3 (
    .in(m2_3),
    .out(m2_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m44_3 (
    .in(m44_3),
    .out(m44_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m28_2 (
    .in(m28_2),
    .out(m28_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m28_3 (
    .in(m28_3),
    .out(m28_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t16_0 (
    .in(t16_0),
    .out(t16_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t16_1 (
    .in(t16_1),
    .out(t16_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t16_2 (
    .in(t16_2),
    .out(t16_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m25_2 (
    .in(m25_2),
    .out(m25_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m25_3 (
    .in(m25_3),
    .out(m25_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m1_1 (
    .in(m1_1),
    .out(m1_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m1_2 (
    .in(m1_2),
    .out(m1_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m1_3 (
    .in(m1_3),
    .out(m1_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m33_3 (
    .in(m33_3),
    .out(m33_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m38_3 (
    .in(m38_3),
    .out(m38_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m15_1 (
    .in(m15_1),
    .out(m15_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m15_2 (
    .in(m15_2),
    .out(m15_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m15_3 (
    .in(m15_3),
    .out(m15_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t15_0 (
    .in(t15_0),
    .out(t15_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t15_1 (
    .in(t15_1),
    .out(t15_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t15_2 (
    .in(t15_2),
    .out(t15_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m14_1 (
    .in(m14_1),
    .out(m14_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m14_2 (
    .in(m14_2),
    .out(m14_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m14_3 (
    .in(m14_3),
    .out(m14_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t25_0 (
    .in(t25_0),
    .out(t25_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m5_1 (
    .in(m5_1),
    .out(m5_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m5_2 (
    .in(m5_2),
    .out(m5_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m5_3 (
    .in(m5_3),
    .out(m5_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t4_0 (
    .in(t4_0),
    .out(t4_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t4_1 (
    .in(t4_1),
    .out(t4_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t4_2 (
    .in(t4_2),
    .out(t4_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m9_1 (
    .in(m9_1),
    .out(m9_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m9_2 (
    .in(m9_2),
    .out(m9_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m9_3 (
    .in(m9_3),
    .out(m9_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m43_3 (
    .in(m43_3),
    .out(m43_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m45_3 (
    .in(m45_3),
    .out(m45_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t17_0 (
    .in(t17_0),
    .out(t17_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t17_1 (
    .in(t17_1),
    .out(t17_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t17_2 (
    .in(t17_2),
    .out(t17_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t1_0 (
    .in(t1_0),
    .out(t1_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t1_1 (
    .in(t1_1),
    .out(t1_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t1_2 (
    .in(t1_2),
    .out(t1_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m27_1 (
    .in(m27_1),
    .out(m27_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m27_2 (
    .in(m27_2),
    .out(m27_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m27_3 (
    .in(m27_3),
    .out(m27_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m8_1 (
    .in(m8_1),
    .out(m8_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m8_2 (
    .in(m8_2),
    .out(m8_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m8_3 (
    .in(m8_3),
    .out(m8_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m11_1 (
    .in(m11_1),
    .out(m11_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m11_2 (
    .in(m11_2),
    .out(m11_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m11_3 (
    .in(m11_3),
    .out(m11_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t10_0 (
    .in(t10_0),
    .out(t10_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t10_1 (
    .in(t10_1),
    .out(t10_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t10_2 (
    .in(t10_2),
    .out(t10_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m24_1 (
    .in(m24_1),
    .out(m24_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m24_2 (
    .in(m24_2),
    .out(m24_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m24_3 (
    .in(m24_3),
    .out(m24_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m21_1 (
    .in(m21_1),
    .out(m21_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m21_2 (
    .in(m21_2),
    .out(m21_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m21_3 (
    .in(m21_3),
    .out(m21_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m42_3 (
    .in(m42_3),
    .out(m42_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m6_1 (
    .in(m6_1),
    .out(m6_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m6_2 (
    .in(m6_2),
    .out(m6_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m6_3 (
    .in(m6_3),
    .out(m6_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t22_0 (
    .in(t22_0),
    .out(t22_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t22_1 (
    .in(t22_1),
    .out(t22_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t22_2 (
    .in(t22_2),
    .out(t22_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m35_3 (
    .in(m35_3),
    .out(m35_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t24_0 (
    .in(t24_0),
    .out(t24_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m41_3 (
    .in(m41_3),
    .out(m41_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m19_1 (
    .in(m19_1),
    .out(m19_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m19_2 (
    .in(m19_2),
    .out(m19_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_m19_3 (
    .in(m19_3),
    .out(m19_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t2_0 (
    .in(t2_0),
    .out(t2_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t2_1 (
    .in(t2_1),
    .out(t2_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_t2_2 (
    .in(t2_2),
    .out(t2_3),
    .clk(clk)
);
endmodule
