`timescale 1ns/1ps

// latency = 4

// Fully pipeline PINI circuit in 4 clock cycles.
// This file has been automatically generated.
`ifdef FULLVERIF
(* fv_prop = "PINI", fv_strat = "composite", fv_order=d *)
`endif
module canright # ( parameter d=2 ) (
    clk,
    i0,
    i1,
    i2,
    i3,
    i4,
    i5,
    i6,
    i7,
    o0,
    o1,
    o2,
    o3,
    o4,
    o5,
    o6,
    o7,
    inverse,
    rnd_0,
    rnd_1,
    rnd_2,
    rnd_3,
);
`include "MSKand_hpc1.vh"
`include "MSKand_hpc2.vh"
`include "MSKand_hpc3.vh"
(* fv_type="clock" *)
input clk;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i0;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i1;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i2;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i3;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i4;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i5;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i6;
(* fv_type="sharing", fv_latency=0, fv_count=1 *)
input [d-1:0] i7;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o0;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o1;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o2;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o3;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o4;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o5;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o6;
(* fv_type="sharing", fv_latency=4, fv_count=1 *)
output [d-1:0] o7;
(* fv_type="random", fv_count=1, fv_rnd_count_0=1*(4*d*(d-1)), fv_rnd_lat_0=0  *)
input [1*(4*d*(d-1))-1:0] rnd_0;
(* fv_type="random", fv_count=1, fv_rnd_count_0=1*(2*d*(d-1)), fv_rnd_lat_0=1  *)
input [1*(2*d*(d-1))-1:0] rnd_1;
(* fv_type="random", fv_count=1, fv_rnd_count_0=2*(2*d*(d-1)), fv_rnd_lat_0=2  *)
input [2*(2*d*(d-1))-1:0] rnd_2;
(* fv_type="random", fv_count=1, fv_rnd_count_0=2*(4*d*(d-1)), fv_rnd_lat_0=3  *)
input [2*(4*d*(d-1))-1:0] rnd_3;
(* fv_type="control", fv_latency=0, fv_count=1 *)
input [1-1:0] inverse;
wire [d-1:0] gen0_0;
wire [d-1:0] gen1_0;
wire [d-1:0] gen10_0;
wire [d-1:0] gen10_1;
wire [d-1:0] gen10_2;
wire [d-1:0] gen10_3;
wire [d-1:0] gen100_4;
wire [d-1:0] gen101_4;
wire [d-1:0] gen102_4;
wire [d-1:0] gen103_4;
wire [d-1:0] gen104_4;
wire [d-1:0] gen105_4;
wire [d-1:0] gen106_4;
wire [d-1:0] gen107_3;
wire [d-1:0] gen107_4;
wire [d-1:0] gen108_3;
wire [d-1:0] gen108_4;
wire [d-1:0] gen109_3;
wire [d-1:0] gen109_4;
wire [d-1:0] gen11_0;
wire [d-1:0] gen110_3;
wire [d-1:0] gen110_4;
wire [d-1:0] gen12_0;
wire [d-1:0] gen13_0;
wire [d-1:0] gen13_1;
wire [d-1:0] gen13_2;
wire [d-1:0] gen13_3;
wire [d-1:0] gen14_0;
wire [d-1:0] gen15_0;
wire [d-1:0] gen16_0;
wire [d-1:0] gen16_1;
wire [d-1:0] gen16_2;
wire [d-1:0] gen16_3;
wire [d-1:0] gen17_0;
wire [d-1:0] gen18_0;
wire [d-1:0] gen19_0;
wire [d-1:0] gen19_1;
wire [d-1:0] gen19_2;
wire [d-1:0] gen19_3;
wire [d-1:0] gen2_0;
wire [d-1:0] gen2_1;
wire [d-1:0] gen2_2;
wire [d-1:0] gen2_3;
wire [d-1:0] gen20_0;
wire [d-1:0] gen21_0;
wire [d-1:0] gen22_0;
wire [d-1:0] gen22_1;
wire [d-1:0] gen22_2;
wire [d-1:0] gen22_3;
wire [d-1:0] gen23_4;
wire [d-1:0] gen24_4;
wire [d-1:0] gen25_4;
wire [d-1:0] gen26_4;
wire [d-1:0] gen27_4;
wire [d-1:0] gen28_4;
wire [d-1:0] gen29_4;
wire [d-1:0] gen3_0;
wire [d-1:0] gen30_4;
wire [d-1:0] gen31_4;
wire [d-1:0] gen32_4;
wire [d-1:0] gen33_4;
wire [d-1:0] gen34_4;
wire [d-1:0] gen35_4;
wire [d-1:0] gen36_4;
wire [d-1:0] gen37_4;
wire [d-1:0] gen38_4;
wire [d-1:0] gen39_4;
wire [d-1:0] gen4_0;
wire [d-1:0] gen40_4;
wire [d-1:0] gen41_4;
wire [d-1:0] gen42_4;
wire [d-1:0] gen43_0;
wire [d-1:0] gen44_0;
wire [d-1:0] gen45_0;
wire [d-1:0] gen46_0;
wire [d-1:0] gen47_0;
wire [d-1:0] gen48_0;
wire [d-1:0] gen49_0;
wire [d-1:0] gen5_0;
wire [d-1:0] gen5_1;
wire [d-1:0] gen5_2;
wire [d-1:0] gen5_3;
wire [d-1:0] gen50_0;
wire [d-1:0] gen51_0;
wire [d-1:0] gen52_0;
wire [d-1:0] gen53_0;
wire [d-1:0] gen54_0;
wire [d-1:0] gen55_0;
wire [d-1:0] gen56_0;
wire [d-1:0] gen57_0;
wire [d-1:0] gen58_0;
wire [d-1:0] gen59_0;
wire [d-1:0] gen6_0;
wire [d-1:0] gen60_0;
wire [d-1:0] gen61_0;
wire [d-1:0] gen62_0;
wire [d-1:0] gen63_0;
wire [d-1:0] gen64_1;
wire [d-1:0] gen64_2;
wire [d-1:0] gen65_1;
wire [d-1:0] gen65_2;
wire [d-1:0] gen66_2;
wire [d-1:0] gen67_1;
wire [d-1:0] gen67_2;
wire [d-1:0] gen68_1;
wire [d-1:0] gen68_2;
wire [d-1:0] gen69_2;
wire [d-1:0] gen7_0;
wire [d-1:0] gen7_1;
wire [d-1:0] gen7_2;
wire [d-1:0] gen7_3;
wire [d-1:0] gen70_2;
wire [d-1:0] gen71_2;
wire [d-1:0] gen72_2;
wire [d-1:0] gen72_3;
wire [d-1:0] gen73_2;
wire [d-1:0] gen74_2;
wire [d-1:0] gen74_3;
wire [d-1:0] gen75_1;
wire [d-1:0] gen76_1;
wire [d-1:0] gen77_1;
wire [d-1:0] gen78_1;
wire [d-1:0] gen79_1;
wire [d-1:0] gen8_0;
wire [d-1:0] gen80_1;
wire [d-1:0] gen81_1;
wire [d-1:0] gen82_1;
wire [d-1:0] gen83_1;
wire [d-1:0] gen84_1;
wire [d-1:0] gen85_1;
wire [d-1:0] gen86_4;
wire [d-1:0] gen87_4;
wire [d-1:0] gen88_4;
wire [d-1:0] gen89_4;
wire [d-1:0] gen9_0;
wire [d-1:0] gen90_4;
wire [d-1:0] gen91_4;
wire [d-1:0] gen92_4;
wire [d-1:0] gen93_4;
wire [d-1:0] gen94_4;
wire [d-1:0] gen95_4;
wire [d-1:0] gen96_4;
wire [d-1:0] gen97_4;
wire [d-1:0] gen98_4;
wire [d-1:0] gen99_4;
wire [d-1:0] i0_0;
wire [d-1:0] i1_0;
wire [d-1:0] i2_0;
wire [d-1:0] i3_0;
wire [d-1:0] i4_0;
wire [d-1:0] i5_0;
wire [d-1:0] i6_0;
wire [d-1:0] i7_0;
wire [d-1:0] o0_4;
wire [d-1:0] o1_4;
wire [d-1:0] o2_4;
wire [d-1:0] o3_4;
wire [d-1:0] o4_4;
wire [d-1:0] o5_4;
wire [d-1:0] o6_4;
wire [d-1:0] o7_4;
assign i0_0 = i0;
assign i1_0 = i1;
assign i2_0 = i2;
assign i3_0 = i3;
assign i4_0 = i4;
assign i5_0 = i5;
assign i6_0 = i6;
assign i7_0 = i7;
assign o0 = o0_4;
assign o1 = o1_4;
assign o2 = o2_4;
assign o3 = o3_4;
assign o4 = o4_4;
assign o5 = o5_4;
assign o6 = o6_4;
assign o7 = o7_4;


wire [1-1:0] inverse_0 = inverse;
reg [1-1:0] inverse_1;
reg [1-1:0] inverse_2;
reg [1-1:0] inverse_3;
reg [1-1:0] inverse_4;
always @(posedge clk) inverse_1 <= inverse_0;
always @(posedge clk) inverse_2 <= inverse_1;
always @(posedge clk) inverse_3 <= inverse_2;
always @(posedge clk) inverse_4 <= inverse_3;


MSKinv #(.d(d)) comp_gen43_0 (
    .out(gen43_0),
    .in(i0_0)
);
MSKinv #(.d(d)) comp_gen44_0 (
    .out(gen44_0),
    .in(i1_0)
);
MSKxor #(.d(d)) comp_gen49_0 (
    .out(gen49_0),
    .ina(i0_0),
    .inb(i1_0)
);
MSKinv #(.d(d)) comp_gen45_0 (
    .out(gen45_0),
    .in(i5_0)
);
MSKxor #(.d(d)) comp_gen53_0 (
    .out(gen53_0),
    .ina(i0_0),
    .inb(i5_0)
);
MSKinv #(.d(d)) comp_gen46_0 (
    .out(gen46_0),
    .in(i6_0)
);
MSKxor #(.d(d)) comp_gen52_0 (
    .out(gen52_0),
    .ina(i0_0),
    .inb(i4_0)
);
MSKxor #(.d(d)) comp_gen21_0 (
    .out(gen21_0),
    .ina(i4_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen58_0 (
    .out(gen58_0),
    .ina(gen43_0),
    .inb(i3_0)
);
MSKxor #(.d(d)) comp_gen59_0 (
    .out(gen59_0),
    .ina(gen43_0),
    .inb(gen44_0)
);
MSKxor #(.d(d)) comp_gen50_0 (
    .out(gen50_0),
    .ina(gen49_0),
    .inb(i3_0)
);
MSKxor #(.d(d)) comp_gen47_0 (
    .out(gen47_0),
    .ina(gen49_0),
    .inb(i2_0)
);
MSKxor #(.d(d)) comp_gen54_0 (
    .out(gen54_0),
    .ina(gen49_0),
    .inb(i5_0)
);
MSKxor #(.d(d)) comp_gen63_0 (
    .out(gen63_0),
    .ina(i2_0),
    .inb(gen45_0)
);
MSKxor #(.d(d)) comp_gen3_0 (
    .out(gen3_0),
    .ina(gen53_0),
    .inb(i6_0)
);
MSKxor #(.d(d)) comp_gen15_0 (
    .out(gen15_0),
    .ina(i4_0),
    .inb(gen46_0)
);
MSKxor #(.d(d)) comp_gen55_0 (
    .out(gen55_0),
    .ina(gen52_0),
    .inb(i5_0)
);
MSKxor #(.d(d)) comp_gen4_0 (
    .out(gen4_0),
    .ina(gen58_0),
    .inb(i4_0)
);
MSKxor #(.d(d)) comp_gen60_0 (
    .out(gen60_0),
    .ina(gen59_0),
    .inb(i3_0)
);
MSKxor #(.d(d)) comp_gen61_0 (
    .out(gen61_0),
    .ina(gen59_0),
    .inb(i4_0)
);
MSKxor #(.d(d)) comp_gen51_0 (
    .out(gen51_0),
    .ina(gen50_0),
    .inb(i4_0)
);
MSKxor #(.d(d)) comp_gen48_0 (
    .out(gen48_0),
    .ina(gen47_0),
    .inb(i3_0)
);
MSKxor #(.d(d)) comp_gen56_0 (
    .out(gen56_0),
    .ina(gen47_0),
    .inb(i5_0)
);
MSKxor #(.d(d)) comp_gen14_0 (
    .out(gen14_0),
    .ina(gen54_0),
    .inb(i6_0)
);
MSKxor #(.d(d)) comp_gen6_0 (
    .out(gen6_0),
    .ina(gen63_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen11_0 (
    .out(gen11_0),
    .ina(gen3_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen9_0 (
    .out(gen9_0),
    .ina(gen15_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen17_0 (
    .out(gen17_0),
    .ina(gen55_0),
    .inb(i6_0)
);
MSKmux #(.d(d)) comp_gen5_0 (
    .out(gen5_0),
    .in_false(gen3_0),
    .in_true(gen4_0),
    .sel(inverse_0)
);
MSKxor #(.d(d)) comp_gen12_0 (
    .out(gen12_0),
    .ina(gen60_0),
    .inb(gen46_0)
);
MSKxor #(.d(d)) comp_gen18_0 (
    .out(gen18_0),
    .ina(gen61_0),
    .inb(gen46_0)
);
MSKxor #(.d(d)) comp_gen62_0 (
    .out(gen62_0),
    .ina(gen61_0),
    .inb(gen45_0)
);
MSKxor #(.d(d)) comp_gen8_0 (
    .out(gen8_0),
    .ina(gen51_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen0_0 (
    .out(gen0_0),
    .ina(gen48_0),
    .inb(i6_0)
);
MSKxor #(.d(d)) comp_gen57_0 (
    .out(gen57_0),
    .ina(gen56_0),
    .inb(i6_0)
);
MSKmux #(.d(d)) comp_gen16_0 (
    .out(gen16_0),
    .in_false(gen14_0),
    .in_true(gen15_0),
    .sel(inverse_0)
);
MSKmux #(.d(d)) comp_gen7_0 (
    .out(gen7_0),
    .in_false(i0_0),
    .in_true(gen6_0),
    .sel(inverse_0)
);
MSKmux #(.d(d)) comp_gen13_0 (
    .out(gen13_0),
    .in_false(gen11_0),
    .in_true(gen12_0),
    .sel(inverse_0)
);
MSKmux #(.d(d)) comp_gen19_0 (
    .out(gen19_0),
    .in_false(gen17_0),
    .in_true(gen18_0),
    .sel(inverse_0)
);
MSKxor #(.d(d)) comp_gen1_0 (
    .out(gen1_0),
    .ina(gen62_0),
    .inb(gen46_0)
);
MSKmux #(.d(d)) comp_gen10_0 (
    .out(gen10_0),
    .in_false(gen8_0),
    .in_true(gen9_0),
    .sel(inverse_0)
);
MSKxor #(.d(d)) comp_gen20_0 (
    .out(gen20_0),
    .ina(gen57_0),
    .inb(i7_0)
);
MSKxor #(.d(d)) comp_gen79_1 (
    .out(gen79_1),
    .ina(gen16_1),
    .inb(gen5_1)
);
MSKg16mul_hpc3 #(.d(d)) comp_gen81_1 (
    .out0(gen81_1),
    .out1(gen83_1),
    .out2(gen84_1),
    .out3(gen85_1),
    .rnd(rnd_0[0 +: 4*d*(d-1)]),
    .ina0(gen13_0),
    .ina0_prev(gen13_1),
    .ina1(gen16_0),
    .ina1_prev(gen16_1),
    .ina2(gen19_0),
    .ina2_prev(gen19_1),
    .ina3(gen22_0),
    .ina3_prev(gen22_1),
    .inb0(gen2_0),
    .inb1(gen5_0),
    .inb2(gen7_0),
    .inb3(gen10_0),
    .clk(clk)
);
MSKxor #(.d(d)) comp_gen75_1 (
    .out(gen75_1),
    .ina(gen19_1),
    .inb(gen7_1)
);
MSKmux #(.d(d)) comp_gen2_0 (
    .out(gen2_0),
    .in_false(gen0_0),
    .in_true(gen1_0),
    .sel(inverse_0)
);
MSKmux #(.d(d)) comp_gen22_0 (
    .out(gen22_0),
    .in_false(gen20_0),
    .in_true(gen21_0),
    .sel(inverse_0)
);
MSKxor #(.d(d)) comp_gen76_1 (
    .out(gen76_1),
    .ina(gen13_1),
    .inb(gen2_1)
);
MSKxor #(.d(d)) comp_gen78_1 (
    .out(gen78_1),
    .ina(gen22_1),
    .inb(gen10_1)
);
MSKxor #(.d(d)) comp_gen77_1 (
    .out(gen77_1),
    .ina(gen75_1),
    .inb(gen76_1)
);
MSKxor #(.d(d)) comp_gen65_1 (
    .out(gen65_1),
    .ina(gen76_1),
    .inb(gen81_1)
);
MSKxor #(.d(d)) comp_gen82_1 (
    .out(gen82_1),
    .ina(gen76_1),
    .inb(gen79_1)
);
MSKxor #(.d(d)) comp_gen80_1 (
    .out(gen80_1),
    .ina(gen78_1),
    .inb(gen79_1)
);
MSKxor #(.d(d)) comp_gen67_1 (
    .out(gen67_1),
    .ina(gen77_1),
    .inb(gen85_1)
);
MSKxor #(.d(d)) comp_gen68_1 (
    .out(gen68_1),
    .ina(gen82_1),
    .inb(gen83_1)
);
MSKxor #(.d(d)) comp_gen64_1 (
    .out(gen64_1),
    .ina(gen80_1),
    .inb(gen84_1)
);
MSKxor #(.d(d)) comp_gen69_2 (
    .out(gen69_2),
    .ina(gen67_2),
    .inb(gen68_2)
);
MSKxor #(.d(d)) comp_gen66_2 (
    .out(gen66_2),
    .ina(gen64_2),
    .inb(gen65_2)
);
MSKg4mul_hpc3 #(.d(d)) comp_gen71_2 (
    .out0(gen71_2),
    .out1(gen73_2),
    .rnd(rnd_1[0 +: 2*d*(d-1)]),
    .ina0(gen64_1),
    .ina0_prev(gen64_2),
    .ina1(gen67_1),
    .ina1_prev(gen67_2),
    .inb0(gen65_1),
    .inb1(gen68_1),
    .clk(clk)
);
MSKxor #(.d(d)) comp_gen70_2 (
    .out(gen70_2),
    .ina(gen66_2),
    .inb(gen69_2)
);
MSKxor #(.d(d)) comp_gen74_2 (
    .out(gen74_2),
    .ina(gen69_2),
    .inb(gen73_2)
);
MSKxor #(.d(d)) comp_gen72_2 (
    .out(gen72_2),
    .ina(gen70_2),
    .inb(gen71_2)
);
MSKg4mul_hpc3 #(.d(d)) comp_gen107_3 (
    .out0(gen107_3),
    .out1(gen108_3),
    .rnd(rnd_2[0 +: 2*d*(d-1)]),
    .ina0(gen74_2),
    .ina0_prev(gen74_3),
    .ina1(gen72_2),
    .ina1_prev(gen72_3),
    .inb0(gen65_2),
    .inb1(gen68_2),
    .clk(clk)
);
MSKg4mul_hpc3 #(.d(d)) comp_gen109_3 (
    .out0(gen109_3),
    .out1(gen110_3),
    .rnd(rnd_2[1*(2*d*(d-1)) +: 2*d*(d-1)]),
    .ina0(gen74_2),
    .ina0_prev(gen74_3),
    .ina1(gen72_2),
    .ina1_prev(gen72_3),
    .inb0(gen64_2),
    .inb1(gen67_2),
    .clk(clk)
);
MSKg16mul_hpc3 #(.d(d)) comp_gen89_4 (
    .out0(gen89_4),
    .out1(gen96_4),
    .out2(gen92_4),
    .out3(gen97_4),
    .rnd(rnd_3[0 +: 4*d*(d-1)]),
    .ina0(gen109_3),
    .ina0_prev(gen109_4),
    .ina1(gen110_3),
    .ina1_prev(gen110_4),
    .ina2(gen107_3),
    .ina2_prev(gen107_4),
    .ina3(gen108_3),
    .ina3_prev(gen108_4),
    .inb0(gen2_3),
    .inb1(gen5_3),
    .inb2(gen7_3),
    .inb3(gen10_3),
    .clk(clk)
);
MSKg16mul_hpc3 #(.d(d)) comp_gen91_4 (
    .out0(gen91_4),
    .out1(gen102_4),
    .out2(gen24_4),
    .out3(gen87_4),
    .rnd(rnd_3[1*(4*d*(d-1)) +: 4*d*(d-1)]),
    .ina0(gen109_3),
    .ina0_prev(gen109_4),
    .ina1(gen110_3),
    .ina1_prev(gen110_4),
    .ina2(gen107_3),
    .ina2_prev(gen107_4),
    .ina3(gen108_3),
    .ina3_prev(gen108_4),
    .inb0(gen13_3),
    .inb1(gen16_3),
    .inb2(gen19_3),
    .inb3(gen22_3),
    .clk(clk)
);
MSKxor #(.d(d)) comp_gen90_4 (
    .out(gen90_4),
    .ina(gen87_4),
    .inb(gen89_4)
);
MSKxor #(.d(d)) comp_gen86_4 (
    .out(gen86_4),
    .ina(gen91_4),
    .inb(gen24_4)
);
MSKxor #(.d(d)) comp_gen41_4 (
    .out(gen41_4),
    .ina(gen91_4),
    .inb(gen92_4)
);
MSKxor #(.d(d)) comp_gen37_4 (
    .out(gen37_4),
    .ina(gen87_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen42_4 (
    .out(gen42_4),
    .ina(gen87_4),
    .inb(gen97_4)
);
MSKxor #(.d(d)) comp_gen38_4 (
    .out(gen38_4),
    .ina(gen102_4),
    .inb(gen89_4)
);
MSKxor #(.d(d)) comp_gen98_4 (
    .out(gen98_4),
    .ina(gen102_4),
    .inb(gen24_4)
);
MSKxor #(.d(d)) comp_gen32_4 (
    .out(gen32_4),
    .ina(gen102_4),
    .inb(gen92_4)
);
MSKxor #(.d(d)) comp_gen100_4 (
    .out(gen100_4),
    .ina(gen91_4),
    .inb(gen102_4)
);
MSKxor #(.d(d)) comp_gen26_4 (
    .out(gen26_4),
    .ina(gen102_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen94_4 (
    .out(gen94_4),
    .ina(gen90_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen88_4 (
    .out(gen88_4),
    .ina(gen86_4),
    .inb(gen87_4)
);
MSKinv #(.d(d)) comp_gen33_4 (
    .out(gen33_4),
    .in(gen41_4)
);
MSKxor #(.d(d)) comp_gen31_4 (
    .out(gen31_4),
    .ina(gen37_4),
    .inb(gen97_4)
);
MSKinv #(.d(d)) comp_gen35_4 (
    .out(gen35_4),
    .in(gen42_4)
);
MSKmux #(.d(d)) comp_o7_4 (
    .out(o7_4),
    .in_false(gen37_4),
    .in_true(gen38_4),
    .sel(inverse_4)
);
MSKxor #(.d(d)) comp_gen39_4 (
    .out(gen39_4),
    .ina(gen38_4),
    .inb(gen92_4)
);
MSKxor #(.d(d)) comp_gen40_4 (
    .out(gen40_4),
    .ina(gen38_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen99_4 (
    .out(gen99_4),
    .ina(gen98_4),
    .inb(gen87_4)
);
MSKxor #(.d(d)) comp_gen101_4 (
    .out(gen101_4),
    .ina(gen100_4),
    .inb(gen87_4)
);
MSKxor #(.d(d)) comp_gen95_4 (
    .out(gen95_4),
    .ina(gen94_4),
    .inb(gen92_4)
);
MSKxor #(.d(d)) comp_gen93_4 (
    .out(gen93_4),
    .ina(gen88_4),
    .inb(gen96_4)
);
MSKmux #(.d(d)) comp_o4_4 (
    .out(o4_4),
    .in_false(gen31_4),
    .in_true(gen32_4),
    .sel(inverse_4)
);
MSKinv #(.d(d)) comp_gen23_4 (
    .out(gen23_4),
    .in(gen39_4)
);
MSKinv #(.d(d)) comp_gen25_4 (
    .out(gen25_4),
    .in(gen40_4)
);
MSKxor #(.d(d)) comp_gen28_4 (
    .out(gen28_4),
    .ina(gen40_4),
    .inb(gen97_4)
);
MSKxor #(.d(d)) comp_gen103_4 (
    .out(gen103_4),
    .ina(gen99_4),
    .inb(gen89_4)
);
MSKxor #(.d(d)) comp_gen105_4 (
    .out(gen105_4),
    .ina(gen101_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen29_4 (
    .out(gen29_4),
    .ina(gen95_4),
    .inb(gen97_4)
);
MSKxor #(.d(d)) comp_gen27_4 (
    .out(gen27_4),
    .ina(gen93_4),
    .inb(gen92_4)
);
MSKmux #(.d(d)) comp_o0_4 (
    .out(o0_4),
    .in_false(gen23_4),
    .in_true(gen24_4),
    .sel(inverse_4)
);
MSKmux #(.d(d)) comp_o1_4 (
    .out(o1_4),
    .in_false(gen25_4),
    .in_true(gen26_4),
    .sel(inverse_4)
);
MSKxor #(.d(d)) comp_gen104_4 (
    .out(gen104_4),
    .ina(gen103_4),
    .inb(gen96_4)
);
MSKxor #(.d(d)) comp_gen106_4 (
    .out(gen106_4),
    .ina(gen105_4),
    .inb(gen92_4)
);
MSKmux #(.d(d)) comp_o2_4 (
    .out(o2_4),
    .in_false(gen27_4),
    .in_true(gen28_4),
    .sel(inverse_4)
);
MSKxor #(.d(d)) comp_gen34_4 (
    .out(gen34_4),
    .ina(gen27_4),
    .inb(gen97_4)
);
MSKxor #(.d(d)) comp_gen30_4 (
    .out(gen30_4),
    .ina(gen104_4),
    .inb(gen92_4)
);
MSKxor #(.d(d)) comp_gen36_4 (
    .out(gen36_4),
    .ina(gen106_4),
    .inb(gen97_4)
);
MSKmux #(.d(d)) comp_o5_4 (
    .out(o5_4),
    .in_false(gen33_4),
    .in_true(gen34_4),
    .sel(inverse_4)
);
MSKmux #(.d(d)) comp_o3_4 (
    .out(o3_4),
    .in_false(gen29_4),
    .in_true(gen30_4),
    .sel(inverse_4)
);
MSKmux #(.d(d)) comp_o6_4 (
    .out(o6_4),
    .in_false(gen35_4),
    .in_true(gen36_4),
    .sel(inverse_4)
);
MSKreg #(.d(d)) reg_gen107_3 (
    .in(gen107_3),
    .out(gen107_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen68_1 (
    .in(gen68_1),
    .out(gen68_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen7_0 (
    .in(gen7_0),
    .out(gen7_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen7_1 (
    .in(gen7_1),
    .out(gen7_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen7_2 (
    .in(gen7_2),
    .out(gen7_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen108_3 (
    .in(gen108_3),
    .out(gen108_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen67_1 (
    .in(gen67_1),
    .out(gen67_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen2_0 (
    .in(gen2_0),
    .out(gen2_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen2_1 (
    .in(gen2_1),
    .out(gen2_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen2_2 (
    .in(gen2_2),
    .out(gen2_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen5_0 (
    .in(gen5_0),
    .out(gen5_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen5_1 (
    .in(gen5_1),
    .out(gen5_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen5_2 (
    .in(gen5_2),
    .out(gen5_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen72_2 (
    .in(gen72_2),
    .out(gen72_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen19_0 (
    .in(gen19_0),
    .out(gen19_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen19_1 (
    .in(gen19_1),
    .out(gen19_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen19_2 (
    .in(gen19_2),
    .out(gen19_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen10_0 (
    .in(gen10_0),
    .out(gen10_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen10_1 (
    .in(gen10_1),
    .out(gen10_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen10_2 (
    .in(gen10_2),
    .out(gen10_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen22_0 (
    .in(gen22_0),
    .out(gen22_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen22_1 (
    .in(gen22_1),
    .out(gen22_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen22_2 (
    .in(gen22_2),
    .out(gen22_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen74_2 (
    .in(gen74_2),
    .out(gen74_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen64_1 (
    .in(gen64_1),
    .out(gen64_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen13_0 (
    .in(gen13_0),
    .out(gen13_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen13_1 (
    .in(gen13_1),
    .out(gen13_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen13_2 (
    .in(gen13_2),
    .out(gen13_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen16_0 (
    .in(gen16_0),
    .out(gen16_1),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen16_1 (
    .in(gen16_1),
    .out(gen16_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen16_2 (
    .in(gen16_2),
    .out(gen16_3),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen109_3 (
    .in(gen109_3),
    .out(gen109_4),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen65_1 (
    .in(gen65_1),
    .out(gen65_2),
    .clk(clk)
);
MSKreg #(.d(d)) reg_gen110_3 (
    .in(gen110_3),
    .out(gen110_4),
    .clk(clk)
);
endmodule
